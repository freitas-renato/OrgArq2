-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
-- CREATED		"Wed Sep 18 19:43:49 2019"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY dataflow IS 
	PORT
	(
		Reg2Loc :  IN  STD_LOGIC;
		branch :  IN  STD_LOGIC;
		memToReg :  IN  STD_LOGIC;
		aluSrc :  IN  STD_LOGIC;
		regWrite :  IN  STD_LOGIC;
		reset :  IN  STD_LOGIC;
		clock :  IN  STD_LOGIC;
		mem_w :  IN  STD_LOGIC;
		mem_r :  IN  STD_LOGIC;
		aluCtl :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		instruction31to21 :  OUT  STD_LOGIC_VECTOR(10 DOWNTO 0)
	);
END dataflow;

ARCHITECTURE bdf_type OF dataflow IS 

COMPONENT estagio_if
	PORT(clock : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 PCSrc : IN STD_LOGIC;
		 Add1Out : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 IMemOut : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PC : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT if_id
	PORT(clock : IN STD_LOGIC;
		 I_IMem : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 I_PC : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_IMem : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 O_PC : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT estagio_id
	PORT(clock : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 Reg2Loc : IN STD_LOGIC;
		 I_regWrite : IN STD_LOGIC;
		 I_instruction4to0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 I_PC : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 instruction : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Mux3Out : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 instruction31to21 : OUT STD_LOGIC_VECTOR(10 DOWNTO 0);
		 O_instruction4to0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 O_PC : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 Reg_Alu : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 Reg_Mux2 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 SEOut : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT id_ex
	PORT(clock : IN STD_LOGIC;
		 I_branch : IN STD_LOGIC;
		 I_mem_w : IN STD_LOGIC;
		 I_mem_r : IN STD_LOGIC;
		 I_memToReg : IN STD_LOGIC;
		 I_aluSrc : IN STD_LOGIC;
		 I_regWrite : IN STD_LOGIC;
		 I_aluCtl : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 I_instruction31to21 : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 I_instruction4to0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 I_PC : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 I_Reg_Alu : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 I_Reg_Mux2 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 I_SEOut : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_branch : OUT STD_LOGIC;
		 O_mem_w : OUT STD_LOGIC;
		 O_mem_r : OUT STD_LOGIC;
		 O_memToReg : OUT STD_LOGIC;
		 O_aluSrc : OUT STD_LOGIC;
		 O_regWrite : OUT STD_LOGIC;
		 O_aluCtl : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 O_instruction31to21 : OUT STD_LOGIC_VECTOR(10 DOWNTO 0);
		 O_instruction4to0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 O_PC : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_Reg_Alu : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_Reg_Mux2 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_SEOut : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT estagio_ex
	PORT(alu_Src : IN STD_LOGIC;
		 I_branch : IN STD_LOGIC;
		 I_mem_w : IN STD_LOGIC;
		 I_mem_r : IN STD_LOGIC;
		 I_memToReg : IN STD_LOGIC;
		 I_regWrite : IN STD_LOGIC;
		 Instruction31to21In : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		 Instruction4to0In : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 PC : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 Reg_Alu : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 Reg_Mux2In : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 SelecaoALU : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 SEOut : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 ZeroAlu : OUT STD_LOGIC;
		 O_branch : OUT STD_LOGIC;
		 O_mem_w : OUT STD_LOGIC;
		 O_mem_r : OUT STD_LOGIC;
		 O_memToReg : OUT STD_LOGIC;
		 O_regWrite : OUT STD_LOGIC;
		 Add1Out : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 AluOut : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 Instruction4to0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 Reg_Mux2 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ex_mem
	PORT(clock : IN STD_LOGIC;
		 I_ZeroAlu : IN STD_LOGIC;
		 I_branch : IN STD_LOGIC;
		 I_mem_w : IN STD_LOGIC;
		 I_mem_r : IN STD_LOGIC;
		 I_memToReg : IN STD_LOGIC;
		 I_regWrite : IN STD_LOGIC;
		 I_Add1 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 I_Alu : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 I_Instruction4to0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 I_Reg_Mux2 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_ZeroAlu : OUT STD_LOGIC;
		 O_branch : OUT STD_LOGIC;
		 O_mem_w : OUT STD_LOGIC;
		 O_mem_r : OUT STD_LOGIC;
		 O_memToReg : OUT STD_LOGIC;
		 O_regWrite : OUT STD_LOGIC;
		 O_Add1 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_Alu : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_Instruction4to0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 O_Reg_Mux2 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT estagio_mem
	PORT(clock : IN STD_LOGIC;
		 mem_w : IN STD_LOGIC;
		 mem_r : IN STD_LOGIC;
		 branch : IN STD_LOGIC;
		 I_RegWrite : IN STD_LOGIC;
		 I_MemToReg : IN STD_LOGIC;
		 ZeroAlu : IN STD_LOGIC;
		 I_Add1Out : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 I_AluOut : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 I_instruction4to0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 Reg_Mux2 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 PC_src : OUT STD_LOGIC;
		 O_MemToReg : OUT STD_LOGIC;
		 O_RegWrite : OUT STD_LOGIC;
		 DMEmOut : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_Add1Out : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_AluOut : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_instruction4to0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mem_wb
	PORT(clock : IN STD_LOGIC;
		 I_RegWrite : IN STD_LOGIC;
		 I_MemToReg : IN STD_LOGIC;
		 I_Alu : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 I_DMEm : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 I_instruction4to0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 O_RegWrite : OUT STD_LOGIC;
		 O_MemToReg : OUT STD_LOGIC;
		 O_Alu : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_DMEm : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 O_instruction4to0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT estagio_wb
	PORT(MemtoReg : IN STD_LOGIC;
		 I_RegWrite : IN STD_LOGIC;
		 AluOut : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 DMemOut : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 Instruction4to0In : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 O_RegWrite : OUT STD_LOGIC;
		 Instruction4to0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 Mux3Out : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC_VECTOR(4 DOWNTO 0);


BEGIN 
instruction31to21 <= SYNTHESIZED_WIRE_9;



b2v_inst : estagio_if
PORT MAP(clock => clock,
		 reset => reset,
		 PCSrc => SYNTHESIZED_WIRE_0,
		 Add1Out => SYNTHESIZED_WIRE_1,
		 IMemOut => SYNTHESIZED_WIRE_2,
		 PC => SYNTHESIZED_WIRE_3);


b2v_inst1 : if_id
PORT MAP(clock => clock,
		 I_IMem => SYNTHESIZED_WIRE_2,
		 I_PC => SYNTHESIZED_WIRE_3,
		 O_IMem => SYNTHESIZED_WIRE_7,
		 O_PC => SYNTHESIZED_WIRE_6);


b2v_inst2 : estagio_id
PORT MAP(clock => clock,
		 reset => reset,
		 Reg2Loc => Reg2Loc,
		 I_regWrite => SYNTHESIZED_WIRE_4,
		 I_instruction4to0 => SYNTHESIZED_WIRE_5,
		 I_PC => SYNTHESIZED_WIRE_6,
		 instruction => SYNTHESIZED_WIRE_7,
		 Mux3Out => SYNTHESIZED_WIRE_8,
		 instruction31to21 => SYNTHESIZED_WIRE_9,
		 O_instruction4to0 => SYNTHESIZED_WIRE_10,
		 O_PC => SYNTHESIZED_WIRE_11,
		 Reg_Alu => SYNTHESIZED_WIRE_12,
		 Reg_Mux2 => SYNTHESIZED_WIRE_13,
		 SEOut => SYNTHESIZED_WIRE_14);


b2v_inst3 : id_ex
PORT MAP(clock => clock,
		 I_branch => branch,
		 I_mem_w => mem_w,
		 I_mem_r => mem_r,
		 I_memToReg => memToReg,
		 I_aluSrc => aluSrc,
		 I_regWrite => regWrite,
		 I_aluCtl => aluCtl,
		 I_instruction31to21 => SYNTHESIZED_WIRE_9,
		 I_instruction4to0 => SYNTHESIZED_WIRE_10,
		 I_PC => SYNTHESIZED_WIRE_11,
		 I_Reg_Alu => SYNTHESIZED_WIRE_12,
		 I_Reg_Mux2 => SYNTHESIZED_WIRE_13,
		 I_SEOut => SYNTHESIZED_WIRE_14,
		 O_branch => SYNTHESIZED_WIRE_16,
		 O_mem_w => SYNTHESIZED_WIRE_17,
		 O_mem_r => SYNTHESIZED_WIRE_18,
		 O_memToReg => SYNTHESIZED_WIRE_19,
		 O_aluSrc => SYNTHESIZED_WIRE_15,
		 O_regWrite => SYNTHESIZED_WIRE_20,
		 O_aluCtl => SYNTHESIZED_WIRE_26,
		 O_instruction31to21 => SYNTHESIZED_WIRE_21,
		 O_instruction4to0 => SYNTHESIZED_WIRE_22,
		 O_PC => SYNTHESIZED_WIRE_23,
		 O_Reg_Alu => SYNTHESIZED_WIRE_24,
		 O_Reg_Mux2 => SYNTHESIZED_WIRE_25,
		 O_SEOut => SYNTHESIZED_WIRE_27);


b2v_inst4 : estagio_ex
PORT MAP(alu_Src => SYNTHESIZED_WIRE_15,
		 I_branch => SYNTHESIZED_WIRE_16,
		 I_mem_w => SYNTHESIZED_WIRE_17,
		 I_mem_r => SYNTHESIZED_WIRE_18,
		 I_memToReg => SYNTHESIZED_WIRE_19,
		 I_regWrite => SYNTHESIZED_WIRE_20,
		 Instruction31to21In => SYNTHESIZED_WIRE_21,
		 Instruction4to0In => SYNTHESIZED_WIRE_22,
		 PC => SYNTHESIZED_WIRE_23,
		 Reg_Alu => SYNTHESIZED_WIRE_24,
		 Reg_Mux2In => SYNTHESIZED_WIRE_25,
		 SelecaoALU => SYNTHESIZED_WIRE_26,
		 SEOut => SYNTHESIZED_WIRE_27,
		 ZeroAlu => SYNTHESIZED_WIRE_28,
		 O_branch => SYNTHESIZED_WIRE_29,
		 O_mem_w => SYNTHESIZED_WIRE_30,
		 O_mem_r => SYNTHESIZED_WIRE_31,
		 O_memToReg => SYNTHESIZED_WIRE_32,
		 O_regWrite => SYNTHESIZED_WIRE_33,
		 Add1Out => SYNTHESIZED_WIRE_34,
		 AluOut => SYNTHESIZED_WIRE_35,
		 Instruction4to0 => SYNTHESIZED_WIRE_36,
		 Reg_Mux2 => SYNTHESIZED_WIRE_37);


b2v_inst5 : ex_mem
PORT MAP(clock => clock,
		 I_ZeroAlu => SYNTHESIZED_WIRE_28,
		 I_branch => SYNTHESIZED_WIRE_29,
		 I_mem_w => SYNTHESIZED_WIRE_30,
		 I_mem_r => SYNTHESIZED_WIRE_31,
		 I_memToReg => SYNTHESIZED_WIRE_32,
		 I_regWrite => SYNTHESIZED_WIRE_33,
		 I_Add1 => SYNTHESIZED_WIRE_34,
		 I_Alu => SYNTHESIZED_WIRE_35,
		 I_Instruction4to0 => SYNTHESIZED_WIRE_36,
		 I_Reg_Mux2 => SYNTHESIZED_WIRE_37,
		 O_ZeroAlu => SYNTHESIZED_WIRE_43,
		 O_branch => SYNTHESIZED_WIRE_40,
		 O_mem_w => SYNTHESIZED_WIRE_38,
		 O_mem_r => SYNTHESIZED_WIRE_39,
		 O_memToReg => SYNTHESIZED_WIRE_42,
		 O_regWrite => SYNTHESIZED_WIRE_41,
		 O_Add1 => SYNTHESIZED_WIRE_44,
		 O_Alu => SYNTHESIZED_WIRE_45,
		 O_Instruction4to0 => SYNTHESIZED_WIRE_46,
		 O_Reg_Mux2 => SYNTHESIZED_WIRE_47);


b2v_inst6 : estagio_mem
PORT MAP(clock => clock,
		 mem_w => SYNTHESIZED_WIRE_38,
		 mem_r => SYNTHESIZED_WIRE_39,
		 branch => SYNTHESIZED_WIRE_40,
		 I_RegWrite => SYNTHESIZED_WIRE_41,
		 I_MemToReg => SYNTHESIZED_WIRE_42,
		 ZeroAlu => SYNTHESIZED_WIRE_43,
		 I_Add1Out => SYNTHESIZED_WIRE_44,
		 I_AluOut => SYNTHESIZED_WIRE_45,
		 I_instruction4to0 => SYNTHESIZED_WIRE_46,
		 Reg_Mux2 => SYNTHESIZED_WIRE_47,
		 PC_src => SYNTHESIZED_WIRE_0,
		 O_MemToReg => SYNTHESIZED_WIRE_49,
		 O_RegWrite => SYNTHESIZED_WIRE_48,
		 DMEmOut => SYNTHESIZED_WIRE_51,
		 O_Add1Out => SYNTHESIZED_WIRE_1,
		 O_AluOut => SYNTHESIZED_WIRE_50,
		 O_instruction4to0 => SYNTHESIZED_WIRE_52);


b2v_inst7 : mem_wb
PORT MAP(clock => clock,
		 I_RegWrite => SYNTHESIZED_WIRE_48,
		 I_MemToReg => SYNTHESIZED_WIRE_49,
		 I_Alu => SYNTHESIZED_WIRE_50,
		 I_DMEm => SYNTHESIZED_WIRE_51,
		 I_instruction4to0 => SYNTHESIZED_WIRE_52,
		 O_RegWrite => SYNTHESIZED_WIRE_54,
		 O_MemToReg => SYNTHESIZED_WIRE_53,
		 O_Alu => SYNTHESIZED_WIRE_55,
		 O_DMEm => SYNTHESIZED_WIRE_56,
		 O_instruction4to0 => SYNTHESIZED_WIRE_57);


b2v_inst8 : estagio_wb
PORT MAP(MemtoReg => SYNTHESIZED_WIRE_53,
		 I_RegWrite => SYNTHESIZED_WIRE_54,
		 AluOut => SYNTHESIZED_WIRE_55,
		 DMemOut => SYNTHESIZED_WIRE_56,
		 Instruction4to0In => SYNTHESIZED_WIRE_57,
		 O_RegWrite => SYNTHESIZED_WIRE_4,
		 Instruction4to0 => SYNTHESIZED_WIRE_5,
		 Mux3Out => SYNTHESIZED_WIRE_8);


END bdf_type;